module sum_binary(
	input wire a,
	input wire b,
	output wire c);
	
	assign c = b+ a;
	
endmodule