library verilog;
use verilog.vl_types.all;
entity sum_tb is
end sum_tb;
