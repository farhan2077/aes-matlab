library verilog;
use verilog.vl_types.all;
entity arithmetic_operators is
end arithmetic_operators;
